

/*
Q14:Write a constraint on two dimensional array for generating even
 numbers in the first 4 locations and odd numbers in the next 4
 locations.Also the even number should be in multiple of 4 and odd number
 should be multiple of 3 ?
*/



// Q15.	Write a constraint to generate an array with unique values and multiples of 3 ?


// Q16.	Write a constraint to generate unique numbers in an array without using the "unique" keyword ?

// Q17.	Write a constraint to generate prime numbers between the range of 1 to 100 ?
// Q18.	Write a constraint to generate a variable with 0-31 bits as 1 and 32-61 bits as 0 ?
// Q19.	Write a constraint to generate consecutive and non-consecutive elements in a fixed-size array ?
// Q20. Write a constraint to randomly generate 10 unique numbers between 99 and 100 ?
// Q21.	Write a constraint such that the array size is between 5 to 10, and the values are in ascending order ?
// Q22.	Write a constraint to generate even numbers between 10 to 30 using a fixed-size array, dynamic array, and queue ?

// 24.	Write a constraint demonstrating the use of the "solve before" constraint ?
// 25.	Write a code to generate unique elements in an array without using the "unique" keyword or constraints ?
// 26.	Write a constraint for a 2D dynamic array to print consecutive elements ?
// 27.	Write a constraint to check whether the randomized number is a palindrome ?
// 28.	Write a constraint to generate the Fibonacci sequence ?
// 29.	Write a code to check whether the randomized number is an Armstrong number ?
// 30.	Write a constraint so that the elements in two queues are different ?
// 31.	Write a constraint for a variable where the range 0-100 is 70% and 101-255 is 30% ?
